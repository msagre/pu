entity cpu4fpga is
  port (
    clk
